module hex_to_7seg (out1, out2, out3, in);

	output [6:0] out1;
	output [6:0] out2;
	output [6:0] out3;
	input [9:0] in;
	
	reg [6:0] out1;
	reg [6:0] out2;
	reg [6:0] out3;
	
	always @ (*)
		case(in)
		
		10'h0: out1 = 7'b1000000;				// -- 0 --
		10'h1: out1 = 7'b1111001;				// │		 │
		10'h2: out1 = 7'b0100100;				// 5	    1
		10'h3: out1 = 7'b0110000;				// │      │
		10'h4: out1 = 7'b0011001;				// -- 6 --
		10'h5: out1 = 7'b0010010;				// │      │
		10'h6: out1 = 7'b0000010;				// 4      2
		10'h7: out1 = 7'b1111000;				// │      │
		10'h8: out1 = 7'b0000000;				// -- 3 --
		10'h9: out1 = 7'b0011000;
		10'ha: out1 = 7'b0001000;
		10'hb: out1 = 7'b0000011;
		10'hc: out1 = 7'b1000110;
		10'hd: out1 = 7'b0100001;
		10'he: out1 = 7'b0000110;
		10'hf: out1 = 7'b0001110;
		
		
		10'h10: out2 = 7'b1000000;				// -- 0 --
		10'h10: out1 = 7'b1111001;
		10'h1: out2 = 7'b1111001;				// │		 │
		10'h2: out2 = 7'b0100100;				// 5	    1
		10'h3: out2 = 7'b0110000;				// │      │
		10'h4: out2 = 7'b0011001;				// -- 6 --
		10'h5: out2 = 7'b0010010;				// │      │
		10'h6: out2 = 7'b0000010;				// 4      2
		10'h7: out2 = 7'b1111000;				// │      │
		10'h8: out2 = 7'b0000000;				// -- 3 --
		10'h9: out2 = 7'b0011000;
		10'ha: out2 = 7'b0001000;
		10'hb: out2 = 7'b0000011;
		10'hc: out2 = 7'b1000110;
		10'hd: out2 = 7'b0100001;
		10'he: out2 = 7'b0000110;
		10'hf: out2 = 7'b0001110;
		
		
		10'h0: out3 = 7'b1000000;				// -- 0 --
		10'h1: out3 = 7'b1111001;				// │		 │
		10'h2: out3 = 7'b0100100;				// 5	    1
		10'h3: out3 = 7'b0110000;				// │      │
		10'h4: out3 = 7'b0011001;				// -- 6 --
		10'h5: out3 = 7'b0010010;				// │      │
		10'h6: out3 = 7'b0000010;				// 4      2
		10'h7: out3 = 7'b1111000;				// │      │
		10'h8: out3 = 7'b0000000;				// -- 3 --
		10'h9: out3 = 7'b0011000;
		10'ha: out3 = 7'b0001000;
		10'hb: out3 = 7'b0000011;
		10'hc: out3 = 7'b1000110;
		10'hd: out3 = 7'b0100001;
		10'he: out3 = 7'b0000110;
		10'hf: out3 = 7'b0001110;
		endcase
		
endmodule
