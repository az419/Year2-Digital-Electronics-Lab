module hex_to_7seg_DP(decimal);
	
	output decimal;
	
	wire decimal;
	assign decimal = 1'b0;

endmodule